module ks1(a, b, d);
    input [0:0] a, b;
    output[0:0] d;

    assign d = a & b;

endmodule